library verilog;
use verilog.vl_types.all;
entity microprocessor_tb is
end microprocessor_tb;
