library verilog;
use verilog.vl_types.all;
entity GeneralDatapath_tb is
end GeneralDatapath_tb;
