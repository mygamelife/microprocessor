library verilog;
use verilog.vl_types.all;
entity RAM_8bits_tb is
end RAM_8bits_tb;
